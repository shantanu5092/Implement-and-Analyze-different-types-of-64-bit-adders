`timescale 1ns/1ps
module cla64b(op1,op2,sum,clock,crout,reset);
input [63:0] op1,op2;
input clock;
input reset;
output reg crout;
output reg [63:0]sum;

wire [63:0] out1,p;
wire out2;
reg [63:0] in1,in2;
wire [62:0] cout;
wire [15:0] G,P;

always @(posedge clock or posedge reset) begin
            if(reset==1) begin
             in1    <= 64'b0;
	     //$display ("op1 = %h", in1);
             in2    <= 64'b0;
	     //$display ("op2 = %h", in2);
             sum   <= 64'b0;
	     //$display ("sum = %h", out1);
             crout <= 1'b0;
	     //$display ("crout = %h", out2);
             end
             else begin
             in1     <= op1;
             $display ("op1 = %h", in1);
             in2     <= op2;
             $display ("op2 = %h", in2);
             sum   <= out1;
             $display ("sum = %h", out1);
             crout <= out2;
             $display ("crout = %h", out2);
             end
        end

cla_gp gp0 (in1[3:0],in2[3:0],G[0],P[0],cout[2:0],p[3:0]);
cla_gpc gp1 (in1[7:4],in2[7:4],cout[3],G[1],P[1],cout[6:4],p[7:4]);
cla_gpc gp2 (in1[11:8],in2[11:8],cout[7],G[2],P[2],cout[10:8],p[11:8]);
cla_gpc gp3 (in1[15:12],in2[15:12],cout[11],G[3],P[3],cout[14:12],p[15:12]);
cla_gpc gp4 (in1[19:16],in2[19:16],cout[15],G[4],P[4],cout[18:16],p[19:16]);
cla_gpc gp5 (in1[23:20],in2[23:20],cout[19],G[5],P[5],cout[22:20],p[23:20]);
cla_gpc gp6 (in1[27:24],in2[27:24],cout[23],G[6],P[6],cout[26:24],p[27:24]);
cla_gpc gp7 (in1[31:28],in2[31:28],cout[27],G[7],P[7],cout[30:28],p[31:28]);
cla_gpc gp8 (in1[35:32],in2[35:32],cout[31],G[8],P[8],cout[34:32],p[35:32]);
cla_gpc gp9 (in1[39:36],in2[39:36],cout[35],G[9],P[9],cout[38:36],p[39:36]);
cla_gpc gp10 (in1[43:40],in2[43:40],cout[39],G[10],P[10],cout[42:40],p[43:40]);
cla_gpc gp11 (in1[47:44],in2[47:44],cout[43],G[11],P[11],cout[46:44],p[47:44]);
cla_gpc gp12 (in1[51:48],in2[51:48],cout[47],G[12],P[12],cout[50:48],p[51:48]);
cla_gpc gp13 (in1[55:52],in2[55:52],cout[51],G[13],P[13],cout[54:52],p[55:52]);
cla_gpc gp14 (in1[59:56],in2[59:56],cout[55],G[14],P[14],cout[58:56],p[59:56]);
cla_gpc gp15 (in1[63:60],in2[63:60],cout[59],G[15],P[15],cout[62:60],p[63:60]);

  assign cout[3]=G[0];
  assign cout[7]=G[1]|(P[1]&G[0]);
  assign cout[11]=G[2]|(P[2]&G[1])|(P[2]&P[1]&G[0]);
  assign cout[15]=G[3]|(P[3]&G[2])|(P[3]&P[2]&G[1])|(P[3]&P[2]&P[1]&G[0]);
  assign cout[19]=G[4]|(P[4]&G[3])|(P[4]&P[3]&G[2])|(P[4]&P[3]&P[2]&G[1])|(P[4]&P[3]&P[2]&P[1]&G[0]);
  assign cout[23]=G[5]|(P[5]&G[4])|(P[5]&P[4]&G[3])|(P[5]&P[4]&P[3]&G[2])|(P[5]&P[4]&P[3]&P[2]&G[1])|(P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);
  assign cout[27]=G[6]|(P[6]&G[5])|(P[6]&P[5]&G[4])|(P[6]&P[5]&P[4]&G[3])|(P[6]&P[5]&P[4]&P[3]&G[2])|(P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);
  assign cout[31]=G[7]|(P[7]&G[6])|(P[7]&P[6]&G[5])|(P[7]&P[6]&P[5]&G[4])|(P[7]&P[6]&P[5]&P[4]&G[3])|(P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);
  assign cout[35]=G[8]|(P[8]&G[7])|(P[8]&P[7]&G[6])|(P[8]&P[7]&P[6]&G[5])|(P[8]&P[7]&P[6]&P[5]&G[4])|(P[8]&P[7]&P[6]&P[5]&P[4]&G[3])|(P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);
  assign cout[39]=G[9]|(P[9]&G[8])|(P[9]&P[8]&G[7])|(P[9]&P[8]&P[7]&G[6])|(P[9]&P[8]&P[7]&P[6]&G[5])|(P[9]&P[8]&P[7]&P[6]&P[5]&G[4])|(P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3])|(P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);
  assign cout[43]=G[10]|(P[10]&G[9])|(P[10]&P[9]&G[8])|(P[10]&P[9]&P[8]&G[7])|(P[10]&P[9]&P[8]&P[7]&G[6])|(P[10]&P[9]&P[8]&P[7]&P[6]&G[5])|(P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4])|(P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3])|(P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|
  (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);
  assign cout[47]=G[11]|(P[11]&G[10])|(P[11]&P[10]&G[9])|(P[11]&P[10]&P[9]&G[8])|(P[11]&P[10]&P[9]&P[8]&G[7])|(P[11]&P[10]&P[9]&P[8]&P[7]&G[6])|(P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5])|(P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4])|(P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3])|(P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|
  (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);
  assign cout[51]=G[12]|(P[12]&G[11])|(P[12]&P[11]&G[10])|(P[12]&P[11]&P[10]&G[9])|(P[12]&P[11]&P[10]&P[9]&G[8])|(P[12]&P[11]&P[10]&P[9]&P[8]&G[7])|(P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6])|(P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5])|(P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4])|(P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3])|
  (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);
  assign cout[55]=G[13]|(P[13]&G[12])|(P[13]&P[12]&G[11])|(P[13]&P[12]&P[11]&G[10])|(P[13]&P[12]&P[11]&P[10]&G[9])|(P[13]&P[12]&P[11]&P[10]&P[9]&G[8])|(P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7])|(P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6])|(P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5])|(P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4])|
  (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3])|(P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);
  assign cout[59]=G[14]|(P[14]&G[13])|(P[14]&P[13]&G[12])|(P[14]&P[13]&P[12]&G[11])|(P[14]&P[13]&P[12]&P[11]&G[10])|(P[14]&P[13]&P[12]&P[11]&P[10]&G[9])|(P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8])|(P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7])|(P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6])|(P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5])|
  (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4])|(P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3])|(P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);
  assign out2=G[15]|(P[15]&G[14])|(P[15]&P[14]&G[13])|(P[15]&P[14]&P[13]&G[12])|(P[15]&P[14]&P[13]&P[12]&G[11])|(P[15]&P[14]&P[13]&P[12]&P[11]&G[10])|(P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9])|(P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8])|(P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7])|(P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6])|
  (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5])|(P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4])|(P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3])|(P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|
  (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);

  cla_sum su [63:0] (p,{cout,1'b0},out1);

endmodule

module cla_gp(a,b,G,P,cout,p);

input [3:0] a,b;
output G,P;
output [3:0]p;

wire [3:0] g,p;
output [2:0] cout;

assign cout[0]=g[0];
assign cout[1]=g[1]|(p[1]&g[0]);
assign cout[2]=g[2]|(p[2]&g[1])|(p[2]&p[1]&g[0]);


assign G=g[3]|(p[3]&g[2])|(p[3]&p[2]&g[1])|(p[3]&p[2]&p[1]&g[0]);
assign P=p[0]&p[1]&p[2]&p[3];

assign g=a&b;
assign p=a^b;

endmodule

module cla_gpc(a,b,cin,G,P,cout,p);

input [3:0] a,b;
input cin;
output G,P;
output [3:0]p;

wire [3:0] g,p;
output [2:0] cout;

assign cout[0]=g[0]|(p[0]&cin);
assign cout[1]=g[1]|(p[1]&g[0])|(p[0]&p[1]&cin);
assign cout[2]=g[2]|(p[2]&g[1])|(p[2]&p[1]&g[0])|(p[2]&p[1]&p[0]&cin);

assign G=g[3]|(p[3]&g[2])|(p[3]&p[2]&g[1])|(p[3]&p[2]&p[1]&g[0]);
assign P=p[0]&p[1]&p[2]&p[3];

assign g=a&b;
assign p=a^b;

endmodule

module cla_sum(a,b,sum);
input a,b;
output sum;

assign sum=a^b;
endmodule



